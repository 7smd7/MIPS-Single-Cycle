module MipsCPU(clock, reset,PCin,PCout,inst,RegDst, RegWrite, ALUSrc, MemtoReg, MemRead, MemWrite, Branch,      ALUOp,      WriteReg,      ReadData1, ReadData2,      Extend32,      ALU_B,      ShiftOut,      ALUCtl,      Zero,      ALUOut,      Add_ALUOut,      AndGateOut,      ReadData,      WriteData_Reg); 