module AndGate(Branch, Zero, AndGateOut);
    input Branch;
    input Zero;
    output reg AndGateOut;
    always @(*) begin
        AndGateOut <= Branch && Zero;
    end
endmodule