
module MIPS (clock, reset);